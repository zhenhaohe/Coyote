/*
 * Copyright (c) 2021, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Redistribution and use in source and binary forms, with or without modification,
 * are permitted provided that the following conditions are met:
 *
 * 1. Redistributions of source code must retain the above copyright notice,
 * this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright notice,
 * this list of conditions and the following disclaimer in the documentation
 * and/or other materials provided with the distribution.
 * 3. Neither the name of the copyright holder nor the names of its contributors
 * may be used to endorse or promote products derived from this software
 * without specific prior written permission.
 *
 * THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
 * ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
 * THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
 * IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,
 * INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
 * PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
 * HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 * OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE,
 * EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
 */
`timescale 1ns / 1ps

`include "axi_macros.svh"
`include "lynx_macros.svh"

import lynxTypes::*;
import bftTypes::*;

/**
 * User logic
 * 
 */
module auth_role_wrapper #( 
  parameter integer NUM_ENGINE = 4,
  parameter integer VERIFICATION = 0
)(
    AXI4S.s                     s_axis,
    metaIntf.s                  s_meta,

    AXI4S.m                     m_axis,
    metaIntf.m                  m_meta,

    AXI4S.s                     s_key,

    // Clock and reset
    input  wire                 aclk,
    input  wire[0:0]            aresetn
);

AXI4S #(.AXI4S_DATA_BITS(AXI_DATA_BITS)) auth_in();
AXI4S #(.AXI4S_DATA_BITS(AXI_DATA_BITS)) auth_out();


bft_packetizer_ip bft_auth_packetizer_inst(
    .ap_clk(aclk),
    .ap_rst_n(aresetn),
    .s_axis_TREADY ( s_axis.tready ),
    .s_axis_TVALID ( s_axis.tvalid ),
    .s_axis_TDATA ( s_axis.tdata ),
    .s_axis_TKEEP ( s_axis.tkeep ),
    .s_axis_TLAST ( s_axis.tlast ),
    .s_axis_TSTRB (0),
    .s_meta_TVALID (s_meta.valid),
    .s_meta_TREADY (s_meta.ready),
    .s_meta_TDATA (s_meta.data),
    .m_axis_TREADY ( auth_in.tready ),
    .m_axis_TVALID ( auth_in.tvalid ),
    .m_axis_TDATA ( auth_in.tdata ),
    .m_axis_TKEEP ( auth_in.tkeep ),
    .m_axis_TLAST ( auth_in.tlast )
);


auth_role #( 
  .NUM_ENGINE(NUM_ENGINE),
  .VERIFICATION(VERIFICATION)
) auth_role
(
    
    .num_engine(NUM_ENGINE),

    .auth_in_tvalid(auth_in.tvalid),
    .auth_in_tlast(auth_in.tlast),
    .auth_in_tready(auth_in.tready),
    .auth_in_tdata(auth_in.tdata),
    .auth_in_tkeep(auth_in.tkeep),

    .auth_out_tvalid(auth_out.tvalid),
    .auth_out_tlast(auth_out.tlast),
    .auth_out_tready(auth_out.tready),
    .auth_out_tdata(auth_out.tdata),
    .auth_out_tkeep(auth_out.tkeep),

    .auth_key_config_in_tvalid(s_key.tvalid),
    .auth_key_config_in_tlast(s_key.tlast),
    .auth_key_config_in_tready(s_key.tready),
    .auth_key_config_in_tdata(s_key.tdata),
    .auth_key_config_in_tkeep(s_key.tkeep),

    // Clock and reset
    .aclk(aclk),
    .aresetn(aresetn)
);

bft_depacketizer_ip bft_auth_depacketizer (
    .ap_clk(aclk),
    .ap_rst_n(aresetn),
    .s_axis_TREADY ( auth_out.tready ),
    .s_axis_TVALID ( auth_out.tvalid ),
    .s_axis_TDATA ( auth_out.tdata ),
    .s_axis_TKEEP ( auth_out.tkeep ),
    .s_axis_TLAST ( auth_out.tlast ),
    .s_axis_TSTRB (0),
    .m_axis_TREADY ( m_axis.tready ),
    .m_axis_TVALID ( m_axis.tvalid ),
    .m_axis_TDATA ( m_axis.tdata ),
    .m_axis_TKEEP ( m_axis.tkeep ),
    .m_axis_TLAST ( m_axis.tlast ),
    .m_meta_TVALID (m_meta.valid),
    .m_meta_TREADY (m_meta.ready),
    .m_meta_TDATA (m_meta.data)
);


endmodule